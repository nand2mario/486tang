// 486Tang - a port of ao486-MiSTer to Tang Console
// nand2mario, 9/2025
module ao486_top (
    input               clk50,
    input               s0,

    output      [7:0]   led,

    output              UART_TXD,
    input               UART_RXD,

    // SDRAM interface  
    inout       [15:0]  IO_sdram_dq,
    output      [12:0]  O_sdram_addr,
    output      [1:0]   O_sdram_ba,
    output      [1:0]   O_sdram_dqm,
    output              O_sdram_clk,
    output              O_sdram_wen_n,
    output              O_sdram_ras_n,
    output              O_sdram_cas_n,
    output              O_sdram_cs_n,

    // VGA output
    output              vga_clk,
    output reg          vga_hs,
    output reg          vga_vs,
    output reg          vga_de,
    output reg    [7:0] vga_r,
    output reg    [7:0] vga_g,
    output reg    [7:0] vga_b,

    // HDMI output
    output              tmds_clk_n,
    output              tmds_clk_p,
    output        [2:0] tmds_d_n,
    output        [2:0] tmds_d_p,

    // DDR3 interface
    output       [14:0] ddr_addr,
    output        [2:0] ddr_bank,
    output              ddr_cs,
    output              ddr_ras,
    output              ddr_cas,
    output              ddr_we,
    output              ddr_ck,
    output              ddr_ck_n,
    output              ddr_cke,
    output              ddr_odt,
    output              ddr_reset_n,
    output        [1:0] ddr_dm,
    inout        [15:0] ddr_dq,
    inout         [1:0] ddr_dqs,
    inout         [1:0] ddr_dqs_n,

    // SD card
    output              sd_clk,
    inout               sd_cmd,
    inout         [3:0] sd_dat,

    // PS/2 keyboard
    input               ps2_kbclk_in,
    input               ps2_kbdat_in,
    output              ps2_kbclk_out,
    output              ps2_kbdat_out
);

wire clk_sys;       // 20Mhz - 30Mhz main clock
wire clk27;         // for framebuffer DDR3 and HDMI
wire clk_vga;       // generated by ao486_to_hdmi, 74.25Mhz (same as 720p pixel clock)
                    // For 1024x768 @ 60Hz, pixel clock is 65Mhz, so 74.25Mhz is fine.
wire clk_sdram_x2;  // SDRAM logic clock, 2x main clock
wire pll_lock_27;

reg reset = 1'b1;
reg [18:0] reset_counter = {19{1'b1}};

always @(posedge clk_sys) begin
    if (reset_counter == 0) begin
//        if (s0 == 1'b0)
            reset <= 1'b0;
    end else begin
        reset_counter <= reset_counter - 1;
    end
end

// Debug signals from system module
wire [2:0] debug_boot_stage;
wire debug_bios_loaded;
wire debug_vga_bios_sig_bad;
wire debug_first_instruction;
wire debug_sd_error;

pll pll(
   .clkin(clk50), 
   .init_clk(clk50),
   .clkout0(clk_sys),         // main clock
   .clkout1(clk_sdram_x2),    // 2x main clock for SDRAM
   .clkout2(O_sdram_clk)      // 315-degree shifted SDRAM clock   
);

pll_vga pll_vga(
    .clkin(clk50),
    .clkout0(clk_vga),
    .init_clk(clk50)
);

pll_27 pll_27(
    .clkin(clk50),
    .clkout0(clk27),
    .init_clk(clk50),
    .lock(pll_lock_27)
);

localparam VGA_FREQ = 60_000_000;
localparam SYS_FREQ = 27_500_000;

// localparam VGA_FREQ = 74_250_000;
// localparam SYS_FREQ = 25_000_000;
// localparam SYS_FREQ = 20_000_000;

// UART <-> PS/2 bridge (keyboard + mouse + framed TX)
wire [7:0] uart_kbd_data;
wire       uart_kbd_we;
wire [7:0] uart_mouse_data;
wire       uart_mouse_we;
wire [7:0] dbg_uart_byte;
wire       dbg_uart_we;
wire [8:0] mouse_host_cmd;
wire       mouse_host_cmd_rd;

wire vga_ce;
assign vga_clk = vga_ce;

wire clk_audio;
wire [4:0] vol_l;
wire [4:0] vol_r;
wire [4:0] vol_cd_l;
wire [4:0] vol_cd_r;
wire [4:0] vol_midi_l;
wire [4:0] vol_midi_r;
wire [4:0] vol_line_l;
wire [4:0] vol_line_r;
wire [1:0] vol_spk;
wire [4:0] vol_en;              
wire sound_fm_mode = 1'b1;      // OPL3
wire sound_cms_en = 1'b0;

wire speaker_out;

wire [15:0] sb_out_l, sb_out_r;
wire [15:0] opl_out_l, opl_out_r;

// nand2mario: maybe we can just use clk_sys for clk_audio...
pll_audio pll_audio(
    .clkin(clk50),
    .clkout0(clk_audio),
    .init_clk(clk50)
);

system #(.SYS_FREQ(SYS_FREQ)) system (
    .clk_sys(clk_sys),
    .reset(reset),
    .clock_rate(SYS_FREQ),
    .clk_sdram_x2(clk_sdram_x2),

    // SDRAM interface
    .sdram_dq(IO_sdram_dq),
    .sdram_a(O_sdram_addr),
    .sdram_ba(O_sdram_ba),
    .sdram_dqm(O_sdram_dqm),
    .sdram_nwe(O_sdram_wen_n),
    .sdram_nras(O_sdram_ras_n),
    .sdram_ncas(O_sdram_cas_n),
    .sdram_ncs(O_sdram_cs_n),
    .sdram_cke(),            // Always enabled
    .refresh_allowed(1'b1),  // Always allow refresh

    .clk_vga(clk_vga),
    .clock_rate_vga(VGA_FREQ),

    .video_ce(vga_ce),      // TODO: clk_vga needs to be >=2x pixel clock for this to work
    .video_r(vga_r),
    .video_g(vga_g),
    .video_b(vga_b),
    .video_hsync(vga_hs),
    .video_vsync(vga_vs),
    .video_blank_n(vga_de),
    
    // SD card
    .sd_clk(sd_clk),
    .sd_cmd(sd_cmd),
    .sd_dat(sd_dat),

    // UART bridge
    .dbg_uart_byte(dbg_uart_byte),
    .dbg_uart_we(dbg_uart_we),

    // Keyboard injection over UART
    .kbd_data(uart_kbd_data),
    .kbd_data_valid(uart_kbd_we),
    .kbd_host_data(),
    .kbd_host_data_clear(1'b0),

    // Mouse injection over UART
    .mouse_data(uart_mouse_data),
    .mouse_data_valid(uart_mouse_we),
    .mouse_host_cmd(mouse_host_cmd),
    .mouse_host_cmd_clear(mouse_host_cmd_rd),

    // Sound
    .clk_audio(clk_audio),
    .sample_sb_l(sb_out_l),
    .sample_sb_r(sb_out_r),
    .sample_opl_l(opl_out_l),
    .sample_opl_r(opl_out_r),
    .sound_fm_mode(sound_fm_mode),
    .sound_cms_en(sound_cms_en),
    .speaker_out(speaker_out),
    .vol_l(vol_l),
    .vol_r(vol_r),
    .vol_cd_l(vol_cd_l),
    .vol_cd_r(vol_cd_r),
    .vol_midi_l(vol_midi_l),
    .vol_midi_r(vol_midi_r),
    .vol_line_l(vol_line_l),
    .vol_line_r(vol_line_r),
    .vol_spk(vol_spk),
    .vol_en(vol_en),

    // Debug outputs for LEDs
    .debug_boot_stage(debug_boot_stage),
    .debug_bios_loaded(debug_bios_loaded),
    .debug_vga_bios_sig_bad(debug_vga_bios_sig_bad),
    .debug_first_instruction(debug_first_instruction),
    .debug_sd_error(debug_sd_error)
);

reg  [16:0] spk_out;

synchronizer speaker_out_sync
(
	.clk(clk_audio),
	.in(speaker_out),
	.out(speaker_out_clk_audio)
);

reg [15:0] out_l, out_r;
reg [16:0] tmp_l, tmp_r;
always @(posedge clk_audio) begin
	tmp_l <= {opl_out_l[15],opl_out_l} + {sb_out_l[15],sb_out_l} + spk_out;
	tmp_r <= {opl_out_r[15],opl_out_r} + {sb_out_r[15],sb_out_r} + spk_out;
	// clamp the output
	out_l <= (^tmp_l[16:15]) ? {tmp_l[16], {15{tmp_l[15]}}} : tmp_l[15:0];
	out_r <= (^tmp_r[16:15]) ? {tmp_r[16], {15{tmp_r[15]}}} : tmp_r[15:0];
end

uart2ps2 #(.CLK_FREQ(SYS_FREQ), .BAUD(115200)) u_uart2ps2 (
    .clk(clk_sys), .resetn(~reset),
    .uart_rx(UART_RXD), .uart_tx(UART_TXD),
    .kbd_data(uart_kbd_data), .kbd_we(uart_kbd_we),
    .mouse_data(uart_mouse_data), .mouse_we(uart_mouse_we),
    .mouse_host_cmd(mouse_host_cmd), .mouse_host_cmd_rd(mouse_host_cmd_rd),
    .dbg_byte(dbg_uart_byte), .dbg_we(dbg_uart_we)
);

// HDMI output
wire init_calib_complete;
ao486_to_hdmi video (       // DDR3-based framebuffer
	.clk27(clk27), 
    .pll_lock_27(pll_lock_27),
    .clk50(clk50),
    .resetn(1'b1), 
    .clk_pixel(), 
    
    .clk_vga(clk_vga), 
    .vga_r(vga_r), 
    .vga_g(vga_g), 
    .vga_b(vga_b), 
    .vga_hs(vga_hs), 
    .vga_vs(vga_vs), 
    .vga_de(vga_de), 
    .vga_ce(vga_ce),

    .sound_left(out_l),
    .sound_right(out_r),

    .ddr_addr(ddr_addr), 
    .ddr_bank(ddr_bank), 
    .ddr_cs(ddr_cs), 
    .ddr_ras(ddr_ras), 
    .ddr_cas(ddr_cas),
    .ddr_we(ddr_we), 
    .ddr_ck(ddr_ck), 
    .ddr_ck_n(ddr_ck_n), 
    .ddr_cke(ddr_cke), 
    .ddr_odt(ddr_odt),
    .ddr_reset_n(ddr_reset_n), 
    .ddr_dm(ddr_dm), 
    .ddr_dq(ddr_dq), 
    .ddr_dqs(ddr_dqs), 
    .ddr_dqs_n(ddr_dqs_n),

	.tmds_clk_n(tmds_clk_n), 
    .tmds_clk_p(tmds_clk_p), 
    .tmds_d_n(tmds_d_n),
	.tmds_d_p(tmds_d_p),

    .ddr_prefetch_delay(0),         // use default prefetch delay
    .init_calib_complete(init_calib_complete)      // 1: ddr3 is ready
);

// Blink generator for LED indicators (different speeds)
reg [23:0] blink_counter;
always @(posedge clk_sys) blink_counter <= blink_counter + 1;

wire blink_fast = blink_counter[20];    // ~12 Hz blink for VGA BIOS signature error
wire blink_slow = blink_counter[23];    // ~1.5 Hz blink for general use

// Keyboard activity indicator: hold LED for a short time after input
reg [23:0] kbd_timer;
always @(posedge clk_sys) begin
    if (reset) begin
        kbd_timer <= 0;
    end else if (uart_kbd_we) begin
        kbd_timer <= 24'h100000;     
    end else if (kbd_timer != 0) begin
        kbd_timer <= kbd_timer - 1;
    end
end
wire keyboard_active = (kbd_timer != 0);

// SD activity indicator: watch sd_cmd/sd_dat bus transitions
reg [23:0] sd_timer;
reg  [4:0] sd_lines_r;
wire [4:0] sd_lines = {sd_cmd, sd_dat};
always @(posedge clk_sys) begin
    if (reset) begin
        sd_timer  <= 0;
        sd_lines_r <= sd_lines;
    end else begin
        if (sd_lines != sd_lines_r) begin
            sd_lines_r <= sd_lines;
            sd_timer <= 24'h7FFFFF;   // shorter hold for SD activity
        end else if (sd_timer != 0) begin
            sd_timer <= sd_timer - 1;
        end
    end
end
wire sd_active = (sd_timer != 0);

// Sound activity indicator: watch Sound Blaster output for activity
reg [23:0] sound_timer;
reg [15:0] out_l_r, out_r_r;
always @(posedge clk_sys) begin
    if (reset) begin
        sound_timer <= 0;
        out_l_r <= 0;
        out_r_r <= 0;
    end else begin
        out_l_r <= out_l;
        out_r_r <= out_r;
        
        // Detect audio activity: any change in Sound Blaster output or non-zero values
        if ((out_l != out_l_r) || (out_r != out_r_r)) begin
            sound_timer <= 24'h7FFFFF;   // hold for sound activity
        end else if (sound_timer != 0) begin
            sound_timer <= sound_timer - 1;
        end
    end
end
wire sound_active = (sound_timer != 0);

// LED assignment:
// LED 0-2: Boot stage (3-bit binary counter) 
// LED 3: Sound activity (Sound Blaster output)
// LED 4: DDR3 calibration complete
// LED 5: Keyboard activity
// LED 6: SD activity; LED 7: video activity
assign led = ~{
    |vga_r,                                             // LED 7: video red activity
    sd_active,                                          // LED 6: SD activity
    keyboard_active,                                    // LED 5: keyboard input activity
    init_calib_complete,                                // LED 4: DDR3 calibration complete
    sound_active,                                       // LED 3: Sound Blaster activity
    debug_boot_stage                                    // LED 0-2: boot stage (3-bit counter)
};

endmodule
